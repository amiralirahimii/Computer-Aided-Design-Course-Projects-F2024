`timescale 1ns/1ns
module testBench();
	reg clk=0,start=0;
	reg [6:0] X,Y,Z;
	wire done;
	mainProccess	mainProccess(.clk(clk),.start(start),.X(X),.Y(Y),.Z(Z),.done(done));
	always #60 clk=~clk;
	initial begin 
		X=7'b0000100;
		Y=7'b1001010;
		Z=7'b1010100;
		#50 start=1;
		#200 start=0;
		#1200000 $stop;
	end
endmodule
